`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:52:32 12/31/2018 
// Design Name: 
// Module Name:    RegisterFile 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RegisterFile(
    input cs,
    input rd,
    input wr,
    input [2:0] rdReg1,
    input [2:0] rdReg2,
    output [15:0] rdData1,
    output [15:0] rdData2,
    input [15:0] wrData,
    input [2:0] wrReg
    );


endmodule
